library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mips_fd is
    generic ( 
    );
    port
    ( 
    );
end entity;

architecture comportamento of mips_fd is

begin

end architecture;